--This library is free software; you can redistribute it and/or
--modify it under the terms of the GNU Lesser General Public
--License as published by the Free Software Foundation; either
--version 2.1 of the License, or (at your option) any later version.

--This library is distributed in the hope that it will be useful,
--but WITHOUT ANY WARRANTY; without even the implied warranty of
--MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
--Lesser General Public License for more details.

--You should have received a copy of the GNU Lesser General Public
--License along with this library; if not, write to the Free Software
--Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA

-- e_mail : j.l.nunez-yanez@byacom.co.uk

---------------------------------
--  ENTITY       = LEVEL1      --
--  version      = 2.0         --
--  last update  = 1/05/00     --
--  author       = Jose Nunez  --
---------------------------------

-- FUNCTION
--  Top level of the hierarchy.
--  This unit does not include a memory interface

--  PIN LIST
--  START        = indicates start of a compress or decompress operation
--  STOP         = forces the end of the current operation
--  COMPRESS     = selects compression mode
--  DECOMPRESS   = selects decompression mode
--  U_BS_IN      = 15 bits maximum block size 32K. size of the block to be compressed
--  C_BS_INOUT   = 16 bits size of the compressed block. compression read the size of the compressed block. decompresssion input the size of the compressed block. buffers stop when is reached. optional system can non-grant the bus to indicate the same. 
--  CLK          = master clock
--  CLEAR 	     = asynchronous reset generated by the csm
--  U_DATAIN     = data to be compressed
--  C_DATAIN     = data to be decompressed
--  U_DATAOUT    = decompressed data
--  C_DATAOUT    = compressed data
--  ADDR_EN      = enable address tri-states
--  CDATA_EN     = enable compressed data tri-state outputs
--  UDATA_EN     = enable uncompressed data tri-state outputs
--  FINISHED     = signal of finished operation
--  COMPRESSING  = compression mode active
--  FLUSHING     = flush active
--  DECOMPRESSING = decompression active

library ieee, std;
use ieee.std_logic_1164.all;
-- use std.textio.all;

entity level1rc is
	port(
		OVERFLOW_CONTROL    : in  std_logic;
		CS                  : in  std_logic;
		RW                  : in  std_logic;
		ADDRESS             : in  std_logic_vector(1 downto 0);
		--===================================================================================
		--	CONTROL : inout std_logic_vector(31 downto 0);
		CONTROL_IN          : in  std_logic_vector(31 downto 0);
		CONTROL_OUT         : out std_logic_vector(31 downto 0);
		--===================================================================================
		CLK                 : in  std_logic;
		CLEAR               : in  std_logic;
		BUS_ACKNOWLEDGE_U   : in  std_logic;
		BUS_ACKNOWLEDGE_C   : in  std_logic;
		WAIT_U              : in  std_logic;
		WAIT_C              : in  std_logic;
		U_DATAIN            : in  std_logic_vector(31 downto 0);
		C_DATAOUT           : out std_logic_vector(31 downto 0);
		C_DATAOUT_TO_DECOMP : out std_logic_vector(31 downto 0); -- to feedback the data to the decompressor
		FINISHED            : out std_logic;
		COMPRESSING         : out std_logic;
		MODE                : out std_logic; -- to active decompression channel in test mode
		FLUSHING            : out std_logic;
		CODING_OVERFLOW     : out std_logic;
		C_DATA_VALID        : out std_logic;
		CRC_OUT             : out std_logic_vector(31 downto 0);
		BUS_REQUEST_U       : out std_logic;
		BUS_REQUEST_C       : out std_logic
	);
end level1rc;

architecture level1_1 of level1rc is

	-- these are  the components that form level1

	component REG_FILE_C
		port(
			DIN             : in  std_logic_vector(31 downto 0);
			ADDRESS         : in  std_logic_vector(1 downto 0);
			C_BS_IN         : in  std_logic_vector(31 downto 0);
			CRC_IN          : in  std_logic_vector(31 downto 0);
			CLEAR_CR        : in  std_logic;
			FINISH          : in  std_logic;
			RW              : in  std_logic;
			ENABLE          : in  std_logic;
			CLEAR           : in  std_logic;
			CLK             : in  std_logic;
			DOUT            : out std_logic_vector(31 downto 0);
			U_BS_OUT        : out std_logic_vector(31 downto 0);
			CRC_OUT         : out std_logic_vector(31 downto 0);
			START_C         : out std_logic;
			STOP            : out std_logic;
			MODE            : out std_logic;
			THRESHOLD_LEVEL : out std_logic_vector(8 downto 0)
		);
	end component;

	component C_BS_COUNTER_C
		port(
			COMPRESS      : in  std_logic;
			CLEAR         : in  std_logic;
			CLEAR_COUNTER : in  std_logic;
			CLK           : in  std_logic;
			ENABLE_C      : in  std_logic;
			C_BS_OUT      : out std_logic_vector(31 downto 0)
		);

	end component;

	component INPUT_BUFFER_32_32
		port(
			OVERFLOW_CONTROL    : in  std_logic;
			FORCE_STOP          : in  std_logic;
			START               : in  std_logic;
			COMP                : in  std_logic;
			STOP                : in  std_logic;
			READ                : in  std_logic;
			WAITN               : in  std_logic;
			DATA_IN_32          : in  std_logic_vector(31 downto 0);
			BUS_ACKNOWLEDGE     : in  std_logic;
			CLEAR               : in  std_logic;
			CLK                 : in  std_logic;
			DATA_OUT_32         : out std_logic_vector(31 downto 0);
			READY               : out std_logic;
			INC_TC              : out std_logic;
			RESET_TOTAL_COUNTER : out std_logic;
			BUS_REQUEST         : out std_logic
		);
	end component;

	component CRC_UNIT_C_32
		port(DIN     : in  std_logic_vector(31 downto 0);
		     ENABLE  : in  std_logic;
		     CLK     : in  std_logic;
		     RESET   : in  std_logic;
		     CLEAR   : in  std_logic;
		     CRC_OUT : out std_logic_vector(31 downto 0)
		    );
	end component;

	component PARSING_UNIT
		port(
			ENABLE         : in  std_logic; -- buffer is ready
			FINISH         : in  std_logic; -- all the data has been processed
			DATA_IN_32     : in  std_logic_vector(31 downto 0);
			CLEAR          : in  std_logic;
			CLK            : in  std_logic;
			READ           : out std_logic;
			FINISH_PARSING : out std_logic;
			START_ENGINE   : out std_logic;
			MASK           : out std_logic_vector(4 downto 0);
			DATA_OUT_32    : out std_logic_vector(31 downto 0)
		);
	end component;

	component CODING_BUFFER_64_32
		port(
			FORCE_STOP         : in  std_logic;
			START              : in  std_logic;
			FINISHED           : in  std_logic;
			OVERFLOW           : in  std_logic;
			SHORT              : in  std_logic;
			WAITN              : in  std_logic;
			DATA_IN_64         : in  std_logic_vector(63 downto 0);
			THRESHOLD_LEVEL    : in  std_logic_vector(8 downto 0);
			BUS_ACKNOWLEDGE    : in  std_logic;
			CLEAR              : in  std_logic;
			CLK                : in  std_logic;
			DATA_OUT_32        : out std_logic_vector(31 downto 0);
			ENABLE_READ        : out std_logic;
			OVERFLOW_DETECTED  : out std_logic;
			UNDERFLOW_DETECTED : out std_logic;
			FLUSHING           : out std_logic;
			DATA_VALID         : out std_logic;
			FINISH             : out std_logic; -- the buffer process
			BUS_REQUEST        : out std_logic
		);
	end component;

	component csm_c_2
		port(
			START_C       : in  std_logic;
			STOP_C        : in  std_logic;
			FINISH_BUFFER : in  std_logic;
			STOP          : in  std_logic;
			FLUSH_END     : in  std_logic;
			CLK           : in  std_logic;
			CLEAR         : in  std_logic;
			COMP          : out std_logic;
			FLUSH         : out std_logic;
			MOVE_ENABLE   : out std_logic;
			RESET         : out std_logic
		);
	end component;

	component BSL_TC_2_C
		port(
			BLOCK_SIZE : in  std_logic_vector(31 downto 0);
			INC        : in  std_logic;
			CLEAR      : in  std_logic;
			RESET      : in  std_logic;
			CLK        : in  std_logic;
			EO_BLOCK   : out std_logic
		);

	end component;

	component level2_4ca

		port(
			CLK         : in  std_logic;
			CLEAR       : in  std_logic;
			RESET       : in  std_logic;
			COMP        : in  std_logic;
			MOVE_ENABLE : in  std_logic;
			FLUSH       : in  std_logic;
			U_DATAIN    : in  std_logic_vector(31 downto 0);
			MASK        : in  std_logic_vector(4 downto 0);
			FLUSH_END   : out std_logic;
			C_DATAOUT   : out std_logic_vector(63 downto 0);
			SHORT       : out std_logic;
			OVERFLOW    : out std_logic
		);
	end component;

	signal READ_INPUT_BUFFER : std_logic;
	signal OVERFLOW_INT      : std_logic;
	signal MOVE_ENABLE       : std_logic;
	signal FLUSH_INT         : std_logic;
	signal COMP_INT          : std_logic;
	signal LOAD_BS           : std_logic;
	signal INC_TC            : std_logic;
	signal RESET             : std_logic;
	signal EO_BLOCK          : std_logic;
	signal STOP_INT          : std_logic;

	signal START_C_INT               : std_logic;
	signal LATCHED_BS                : std_logic_vector(31 downto 0);
	signal FLUSH_END                 : std_logic;
	signal C_DATAOUT_INT             : std_logic_vector(63 downto 0);
	signal C_DATAOUT_32_INT          : std_logic_vector(31 downto 0);
	signal OVERFLOW_DETECTED_CODING  : std_logic;
	signal UNDERFLOW_DETECTED_CODING : std_logic;
	signal ENABLE_READ               : std_logic;

	signal INC_TC_CSM : std_logic;

	signal BUS_REQUEST_CODING : std_logic;
	signal THRESHOLD_LEVEL    : std_logic_vector(8 downto 0);
	signal FLUSHING_INT       : std_logic;

	signal C_DATA_VALID_INT       : std_logic;
	signal FINISHED_BUFFER_CODING : std_logic;
	signal FINISHED_AUX           : std_logic;
	signal C_BS_OUT               : std_logic_vector(31 downto 0);
	signal CONTROL_AUX            : std_logic_vector(31 downto 0);

	signal PARSER_DATA_IN : std_logic_vector(31 downto 0);

	signal PARSER_DATA_OUT : std_logic_vector(31 downto 0);

	signal MASK : std_logic_vector(4 downto 0);

	signal I_BUFFER_READY      : std_logic;
	signal RESET_TOTAL_COUNTER : std_logic; -- the whole block is reset only once

	signal FINISH_PARSING : std_logic;  -- the parser has parsed all the data

	signal CRC_CODE : std_logic_vector(31 downto 0); -- test mode

	signal START_ENGINE : std_logic;    -- the parser unit starts the engine

	signal SHORT : std_logic;           -- the last output from the compression engine is less or equal to 32 bits

begin

	P_U : PARSING_UNIT
		port map(
			ENABLE         => I_BUFFER_READY,
			FINISH         => RESET_TOTAL_COUNTER, -- all the data has been read from the buffer
			DATA_IN_32     => PARSER_DATA_IN,
			CLEAR          => CLEAR,
			CLK            => CLK,
			READ           => READ_INPUT_BUFFER,
			FINISH_PARSING => FINISH_PARSING,
			START_ENGINE   => START_ENGINE,
			MASK           => MASK,
			DATA_OUT_32    => PARSER_DATA_OUT
		);

	I_B : INPUT_BUFFER_32_32
		port map(
			OVERFLOW_CONTROL    => OVERFLOW_CONTROL,
			FORCE_STOP          => STOP_INT,
			START               => START_C_INT,
			COMP                => COMP_INT,
			STOP                => EO_BLOCK,
			READ                => READ_INPUT_BUFFER,
			WAITN               => WAIT_U,
			DATA_IN_32          => U_DATAIN,
			BUS_ACKNOWLEDGE     => BUS_ACKNOWLEDGE_U,
			CLEAR               => CLEAR,
			CLK                 => CLK,
			DATA_OUT_32         => PARSER_DATA_IN,
			READY               => I_BUFFER_READY,
			INC_TC              => INC_TC,
			RESET_TOTAL_COUNTER => RESET_TOTAL_COUNTER,
			BUS_REQUEST         => BUS_REQUEST_U
		);

	CRC_UNIT_1 : CRC_UNIT_C_32
		port map(DIN     => U_DATAIN,
		         ENABLE  => INC_TC,
		         CLK     => CLK,
		         RESET   => FINISHED_AUX,
		         CLEAR   => CLEAR,
		         CRC_OUT => CRC_CODE
		        );

	level2_4_1 : level2_4ca
		port map(CLK         => CLK,
		         RESET       => RESET,
		         CLEAR       => CLEAR,
		         COMP        => COMP_INT,
		         MOVE_ENABLE => MOVE_ENABLE,
		         FLUSH       => FLUSH_INT,
		         FLUSH_END   => FLUSH_END,
		         MASK        => MASK,
		         C_DATAOUT   => C_DATAOUT_INT,
		         U_DATAIN    => PARSER_DATA_OUT,
		         SHORT       => SHORT,
		         OVERFLOW    => OVERFLOW_INT
		        );

	csm_1 : csm_c_2
		port map(
			START_C       => START_ENGINE,
			STOP_C        => FINISH_PARSING,
			FINISH_BUFFER => RESET_TOTAL_COUNTER,
			STOP          => STOP_INT,
			FLUSH_END     => FLUSH_END,
			CLK           => CLK,
			CLEAR         => CLEAR,
			COMP          => COMP_INT,
			FLUSH         => FLUSH_INT,
			MOVE_ENABLE   => MOVE_ENABLE,
			RESET         => RESET
		);

		-- if decoding underflow active do not increment the counter

	BSL_TC_1 : BSL_TC_2_C
		port map(
			BLOCK_SIZE => LATCHED_BS,
			INC        => INC_TC,
			CLEAR      => CLEAR,
			RESET      => RESET_TOTAL_COUNTER,
			CLK        => CLK,
			EO_BLOCK   => EO_BLOCK
		);

	REG_FILE_1 : REG_FILE_C
		port map(
			DIN             => CONTROL_AUX,
			ADDRESS         => ADDRESS,
			CLEAR_CR        => EO_BLOCK, -- reset the comand register to avoid restart.
			RW              => RW,
			C_BS_IN         => C_BS_OUT,
			CRC_IN          => CRC_CODE,
			FINISH          => FINISHED_BUFFER_CODING,
			ENABLE          => CS,
			CLEAR           => CLEAR,
			CLK             => CLK,
			DOUT            => CONTROL_OUT,
			U_BS_OUT        => LATCHED_BS,
			CRC_OUT         => CRC_OUT,
			START_C         => START_C_INT,
			STOP            => STOP_INT,
			MODE            => MODE,
			THRESHOLD_LEVEL => THRESHOLD_LEVEL
		);

	C_BS_COUNTER_1 : C_BS_COUNTER_C
		port map(
			COMPRESS      => START_C_INT,
			CLEAR_COUNTER => FINISHED_AUX,
			CLEAR         => CLEAR,
			CLK           => CLK,
			ENABLE_C      => C_DATA_VALID_INT,
			C_BS_OUT      => C_BS_OUT
		);

	CODING_BUFFER : CODING_BUFFER_64_32
		port map(
			FORCE_STOP         => STOP_INT,
			START              => COMP_INT,
			FINISHED           => FLUSH_END,
			OVERFLOW           => OVERFLOW_INT,
			SHORT              => SHORT,
			WAITN              => WAIT_C,
			DATA_IN_64         => C_DATAOUT_INT,
			THRESHOLD_LEVEL    => THRESHOLD_LEVEL,
			BUS_ACKNOWLEDGE    => BUS_ACKNOWLEDGE_C,
			CLEAR              => CLEAR,
			CLK                => CLK,
			DATA_OUT_32        => C_DATAOUT_32_INT,
			ENABLE_READ        => ENABLE_READ,
			OVERFLOW_DETECTED  => OVERFLOW_DETECTED_CODING,
			UNDERFLOW_DETECTED => UNDERFLOW_DETECTED_CODING,
			FLUSHING           => FLUSHING_INT,
			FINISH             => FINISHED_BUFFER_CODING,
			DATA_VALID         => C_DATA_VALID_INT,
			BUS_REQUEST        => BUS_REQUEST_CODING
		);

		-- Careful I change this for the PCI implementation
		-- C_DATAOUT <= C_DATAOUT_32_INT when BUS_ACKNOWLEDGE_C = '0' else "ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ";
	C_DATAOUT           <= C_DATAOUT_32_INT;
	C_DATAOUT_TO_DECOMP <= C_DATAOUT_32_INT;
	COMPRESSING         <= COMP_INT;
	FLUSHING            <= FLUSHING_INT;
	BUS_REQUEST_C       <= BUS_REQUEST_CODING;
	FINISHED_AUX        <= FINISHED_BUFFER_CODING;

	C_DATA_VALID <= C_DATA_VALID_INT;

	CODING_OVERFLOW <= OVERFLOW_DETECTED_CODING;

	CONTROL_AUX <= (CONTROL_IN);
	FINISHED    <= FINISHED_AUX;

end level1_1;
